library verilog;
use verilog.vl_types.all;
entity IF_ID is
    port(
        clk_i           : in     vl_logic;
        IR_i            : in     vl_logic_vector(31 downto 0);
        IR_o            : out    vl_logic_vector(31 downto 0);
        isstall_i       : in     vl_logic
    );
end IF_ID;
